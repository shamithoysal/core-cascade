`default_nettype none
`timescale 1ns/1ns

module controller #(
    parameter ADDR_BITS = 8,
    parameter DATA_BITS = 16,
    parameter NUM_CONSUMERS = 4,
    parameter NUM_CHANNELS = 1,
    parameter WRITE_ENABLE = 1
)(
    input  wire clk,
    input  wire reset,

    input  wire [NUM_CONSUMERS-1:0] consumer_read_valid,
    input  wire [ADDR_BITS-1:0] consumer_read_address [NUM_CONSUMERS-1:0],
    output reg  [NUM_CONSUMERS-1:0] consumer_read_ready,
    output reg  [DATA_BITS-1:0] consumer_read_data [NUM_CONSUMERS-1:0],

    input  wire [NUM_CONSUMERS-1:0] consumer_write_valid,
    input  wire [ADDR_BITS-1:0] consumer_write_address [NUM_CONSUMERS-1:0],
    input  wire [DATA_BITS-1:0] consumer_write_data [NUM_CONSUMERS-1:0],
    output reg  [NUM_CONSUMERS-1:0] consumer_write_ready,

    output reg  [NUM_CHANNELS-1:0] mem_read_valid,
    output reg  [ADDR_BITS-1:0] mem_read_address [NUM_CHANNELS-1:0],
    input  wire [NUM_CHANNELS-1:0] mem_read_ready,
    input  wire [DATA_BITS-1:0] mem_read_data [NUM_CHANNELS-1:0],

    output reg  [NUM_CHANNELS-1:0] mem_write_valid,
    output reg  [ADDR_BITS-1:0] mem_write_address [NUM_CHANNELS-1:0],
    output reg  [DATA_BITS-1:0] mem_write_data [NUM_CHANNELS-1:0],
    input  wire [NUM_CHANNELS-1:0] mem_write_ready
);

    localparam IDLE           = 3'b000;
    localparam READ_WAITING   = 3'b010;
    localparam WRITE_WAITING  = 3'b011;
    localparam READ_RELAYING  = 3'b100;
    localparam WRITE_RELAYING = 3'b101;

    reg [2:0] controller_state [NUM_CHANNELS-1:0];
    reg [$clog2(NUM_CONSUMERS)-1:0] current_consumer [NUM_CHANNELS-1:0];
    reg [NUM_CONSUMERS-1:0] channel_serving_consumer;

    integer i, j;

    always @(posedge clk) begin
        if (reset) begin

            mem_read_valid       <= '0;
            mem_write_valid      <= '0;
            consumer_read_ready  <= '0;
            consumer_write_ready <= '0;
            channel_serving_consumer <= '0;

            for (i = 0; i < NUM_CHANNELS; i = i + 1) begin
                mem_read_address[i]  <= '0;
                mem_write_address[i] <= '0;
                mem_write_data[i]    <= '0;
                current_consumer[i]  <= '0;
                controller_state[i]  <= IDLE;
            end

            for (j = 0; j < NUM_CONSUMERS; j = j + 1) begin
                consumer_read_data[j] <= '0;
            end
        end
        else begin

            for (i = 0; i < NUM_CHANNELS; i = i + 1) begin

                case (controller_state[i])

                    IDLE: begin
                        reg found;
                        found = 0;

                        for (j = 0; j < NUM_CONSUMERS; j = j + 1) begin
                            if (!found) begin

                                if (consumer_read_valid[j] &&
                                   !channel_serving_consumer[j]) begin

                                    channel_serving_consumer[j] <= 1'b1;
                                    current_consumer[i]         <= j;

                                    mem_read_valid[i]           <= 1'b1;
                                    mem_read_address[i]         <= consumer_read_address[j];
                                    controller_state[i]         <= READ_WAITING;

                                    found = 1;
                                end
                                else if (WRITE_ENABLE &&
                                         consumer_write_valid[j] &&
                                        !channel_serving_consumer[j]) begin

                                    channel_serving_consumer[j] <= 1'b1;
                                    current_consumer[i]         <= j;

                                    mem_write_valid[i]          <= 1'b1;
                                    mem_write_address[i]        <= consumer_write_address[j];
                                    mem_write_data[i]           <= consumer_write_data[j];
                                    controller_state[i]         <= WRITE_WAITING;

                                    found = 1;
                                end
                            end
                        end
                    end

                    READ_WAITING: begin
                        if (mem_read_ready[i]) begin
                            mem_read_valid[i] <= 1'b0;
                            consumer_read_ready[current_consumer[i]] <= 1'b1;
                            consumer_read_data[current_consumer[i]]  <= mem_read_data[i];
                            controller_state[i] <= READ_RELAYING;
                        end
                    end

                    WRITE_WAITING: begin
                        if (mem_write_ready[i]) begin
                            mem_write_valid[i] <= 1'b0;
                            consumer_write_ready[current_consumer[i]] <= 1'b1;
                            controller_state[i] <= WRITE_RELAYING;
                        end
                    end

                    READ_RELAYING: begin
                        if (!consumer_read_valid[current_consumer[i]]) begin
                            channel_serving_consumer[current_consumer[i]] <= 1'b0;
                            consumer_read_ready[current_consumer[i]] <= 1'b0;
                            controller_state[i] <= IDLE;
                        end
                    end

                    WRITE_RELAYING: begin
                        if (!consumer_write_valid[current_consumer[i]]) begin
                            channel_serving_consumer[current_consumer[i]] <= 1'b0;
                            consumer_write_ready[current_consumer[i]] <= 1'b0;
                            controller_state[i] <= IDLE;
                        end
                    end

                endcase
            end
        end
    end

endmodule
